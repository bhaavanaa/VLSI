// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383
// NAND4 13
// AND3 12
// NAND2 60
// NAND3 14
// AND2 105
// OR2 29
// NOT1 63
// NOR2 61
// BUFF1 26

module c880 (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
             N865,N866,N874,N878,N879,N880);

input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;

output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877;

nand NAND4_1 (N269, N1, N8, N13, N17);
nand NAND4_2 (N270, N1, N26, N13, N17);
and AND3_3 (N273, N29, N36, N42);
and AND3_4 (N276, N1, N26, N51);
nand NAND4_5 (N279, N1, N8, N51, N17);
nand NAND4_6 (N280, N1, N8, N13, N55);
nand NAND4_7 (N284, N59, N42, N68, N72);
nand NAND2_8 (N285, N29, N68);
nand NAND3_9 (N286, N59, N68, N74);
and AND3_10 (N287, N29, N75, N80);
and AND3_11 (N290, N29, N75, N42);
and AND3_12 (N291, N29, N36, N80);
and AND3_13 (N292, N29, N36, N42);
and AND3_14 (N293, N59, N75, N80);
and AND3_15 (N294, N59, N75, N42);
and AND3_16 (N295, N59, N36, N80);
and AND3_17 (N296, N59, N36, N42);
and AND2_18 (N297, N85, N86);
or OR2_19 (N298, N87, N88);
nand NAND2_20 (N301, N91, N96);
or OR2_21 (N302, N91, N96);
nand NAND2_22 (N303, N101, N106);
or OR2_23 (N304, N101, N106);
nand NAND2_24 (N305, N111, N116);
or OR2_25 (N306, N111, N116);
nand NAND2_26 (N307, N121, N126);
or OR2_27 (N308, N121, N126);
and AND2_28 (N309, N8, N138);
not NOT1_29 (N310, N268);
and AND2_30 (N316, N51, N138);
and AND2_31 (N317, N17, N138);
and AND2_32 (N318, N152, N138);
nand NAND2_33 (N319, N59, N156);
nor NOR2_34 (N322, N17, N42);
and AND2_35 (N323, N17, N42);
nand NAND2_36 (N324, N159, N165);
or OR2_37 (N325, N159, N165);
nand NAND2_38 (N326, N171, N177);
or OR2_39 (N327, N171, N177);
nand NAND2_40 (N328, N183, N189);
or OR2_41 (N329, N183, N189);
nand NAND2_42 (N330, N195, N201);
or OR2_43 (N331, N195, N201);
and AND2_44 (N332, N210, N91);
and AND2_45 (N333, N210, N96);
and AND2_46 (N334, N210, N101);
and AND2_47 (N335, N210, N106);
and AND2_48 (N336, N210, N111);
and AND2_49 (N337, N255, N259);
and AND2_50 (N338, N210, N116);
and AND2_51 (N339, N255, N260);
and AND2_52 (N340, N210, N121);
and AND2_53 (N341, N255, N267);
not NOT1_54 (N342, N269);
not NOT1_55 (N343, N273);
or OR2_56 (N344, N270, N273);
not NOT1_57 (N345, N276);
not NOT1_58 (N346, N276);
not NOT1_59 (N347, N279);
nor NOR2_60 (N348, N280, N284);
or OR2_61 (N349, N280, N285);
or OR2_62 (N350, N280, N286);
not NOT1_63 (N351, N293);
not NOT1_64 (N352, N294);
not NOT1_65 (N353, N295);
not NOT1_66 (N354, N296);
nand NAND2_67 (N355, N89, N298);
and AND2_68 (N356, N90, N298);
nand NAND2_69 (N357, N301, N302);
nand NAND2_70 (N360, N303, N304);
nand NAND2_71 (N363, N305, N306);
nand NAND2_72 (N366, N307, N308);
not NOT1_73 (N369, N310);
nor NOR2_74 (N375, N322, N323);
nand NAND2_75 (N376, N324, N325);
nand NAND2_76 (N379, N326, N327);
nand NAND2_77 (N382, N328, N329);
nand NAND2_78 (N385, N330, N331);
buf BUFF1_79 (N388, N290);
buf BUFF1_80 (N389, N291);
buf BUFF1_81 (N390, N292);
buf BUFF1_82 (N391, N297);
or OR2_83 (N392, N270, N343);
not NOT1_84 (N393, N345);
not NOT1_85 (N399, N346);
and AND2_86 (N400, N348, N73);
not NOT1_87 (N401, N349);
not NOT1_88 (N402, N350);
not NOT1_89 (N403, N355);
not NOT1_90 (N404, N357);
not NOT1_91 (N405, N360);
and AND2_92 (N406, N357, N360);
not NOT1_93 (N407, N363);
not NOT1_94 (N408, N366);
and AND2_95 (N409, N363, N366);
nand NAND2_96 (N410, N347, N352);
not NOT1_97 (N411, N376);
not NOT1_98 (N412, N379);
and AND2_99 (N413, N376, N379);
not NOT1_100 (N414, N382);
not NOT1_101 (N415, N385);
and AND2_102 (N416, N382, N385);
and AND2_103 (N417, N210, N369);
buf BUFF1_104 (N418, N342);
buf BUFF1_105 (N419, N344);
buf BUFF1_106 (N420, N351);
buf BUFF1_107 (N421, N353);
buf BUFF1_108 (N422, N354);
buf BUFF1_109 (N423, N356);
not NOT1_110 (N424, N400);
and AND2_111 (N425, N404, N405);
and AND2_112 (N426, N407, N408);
and AND3_113 (N427, N319, N393, N55);
and AND3_114 (N432, N393, N17, N287);
nand NAND3_115 (N437, N393, N287, N55);
nand NAND4_116 (N442, N375, N59, N156, N393);
nand NAND3_117 (N443, N393, N319, N17);
and AND2_118 (N444, N411, N412);
and AND2_119 (N445, N414, N415);
buf BUFF1_120 (N446, N392);
buf BUFF1_121 (N447, N399);
buf BUFF1_122 (N448, N401);
buf BUFF1_123 (N449, N402);
buf BUFF1_124 (N450, N403);
not NOT1_125 (N451, N424);
nor NOR2_126 (N460, N406, N425);
nor NOR2_127 (N463, N409, N426);
nand NAND2_128 (N466, N442, N410);
and AND2_129 (N475, N143, N427);
and AND2_130 (N476, N310, N432);
and AND2_131 (N477, N146, N427);
and AND2_132 (N478, N310, N432);
and AND2_133 (N479, N149, N427);
and AND2_134 (N480, N310, N432);
and AND2_135 (N481, N153, N427);
and AND2_136 (N482, N310, N432);
nand NAND2_137 (N483, N443, N1);
or OR2_138 (N488, N369, N437);
or OR2_139 (N489, N369, N437);
or OR2_140 (N490, N369, N437);
or OR2_141 (N491, N369, N437);
nor NOR2_142 (N492, N413, N444);
nor NOR2_143 (N495, N416, N445);
nand NAND2_144 (N498, N130, N460);
or OR2_145 (N499, N130, N460);
nand NAND2_146 (N500, N463, N135);
or OR2_147 (N501, N463, N135);
and AND2_148 (N502, N91, N466);
nor NOR2_149 (N503, N475, N476);
and AND2_150 (N504, N96, N466);
nor NOR2_151 (N505, N477, N478);
and AND2_152 (N506, N101, N466);
nor NOR2_153 (N507, N479, N480);
and AND2_154 (N508, N106, N466);
nor NOR2_155 (N509, N481, N482);
and AND2_156 (N510, N143, N483);
and AND2_157 (N511, N111, N466);
and AND2_158 (N512, N146, N483);
and AND2_159 (N513, N116, N466);
and AND2_160 (N514, N149, N483);
and AND2_161 (N515, N121, N466);
and AND2_162 (N516, N153, N483);
and AND2_163 (N517, N126, N466);
nand NAND2_164 (N518, N130, N492);
or OR2_165 (N519, N130, N492);
nand NAND2_166 (N520, N495, N207);
or OR2_167 (N521, N495, N207);
and AND2_168 (N522, N451, N159);
and AND2_169 (N523, N451, N165);
and AND2_170 (N524, N451, N171);
and AND2_171 (N525, N451, N177);
and AND2_172 (N526, N451, N183);
nand NAND2_173 (N527, N451, N189);
nand NAND2_174 (N528, N451, N195);
nand NAND2_175 (N529, N451, N201);
nand NAND2_176 (N530, N498, N499);
nand NAND2_177 (N533, N500, N501);
nor NOR2_178 (N536, N309, N502);
nor NOR2_179 (N537, N316, N504);
nor NOR2_180 (N538, N317, N506);
nor NOR2_181 (N539, N318, N508);
nor NOR2_182 (N540, N510, N511);
nor NOR2_183 (N541, N512, N513);
nor NOR2_184 (N542, N514, N515);
nor NOR2_185 (N543, N516, N517);
nand NAND2_186 (N544, N518, N519);
nand NAND2_187 (N547, N520, N521);
not NOT1_188 (N550, N530);
not NOT1_189 (N551, N533);
and AND2_190 (N552, N530, N533);
nand NAND2_191 (N553, N536, N503);
nand NAND2_192 (N557, N537, N505);
nand NAND2_193 (N561, N538, N507);
nand NAND2_194 (N565, N539, N509);
nand NAND2_195 (N569, N488, N540);
nand NAND2_196 (N573, N489, N541);
nand NAND2_197 (N577, N490, N542);
nand NAND2_198 (N581, N491, N543);
not NOT1_199 (N585, N544);
not NOT1_200 (N586, N547);
and AND2_201 (N587, N544, N547);
and AND2_202 (N588, N550, N551);
and AND2_203 (N589, N585, N586);
nand NAND2_204 (N590, N553, N159);
or OR2_205 (N593, N553, N159);
and AND2_206 (N596, N246, N553);
nand NAND2_207 (N597, N557, N165);
or OR2_208 (N600, N557, N165);
and AND2_209 (N605, N246, N557);
nand NAND2_210 (N606, N561, N171);
or OR2_211 (N609, N561, N171);
and AND2_212 (N615, N246, N561);
nand NAND2_213 (N616, N565, N177);
or OR2_214 (N619, N565, N177);
and AND2_215 (N624, N246, N565);
nand NAND2_216 (N625, N569, N183);
or OR2_217 (N628, N569, N183);
and AND2_218 (N631, N246, N569);
nand NAND2_219 (N632, N573, N189);
or OR2_220 (N635, N573, N189);
and AND2_221 (N640, N246, N573);
nand NAND2_222 (N641, N577, N195);
or OR2_223 (N644, N577, N195);
and AND2_224 (N650, N246, N577);
nand NAND2_225 (N651, N581, N201);
or OR2_226 (N654, N581, N201);
and AND2_227 (N659, N246, N581);
nor NOR2_228 (N660, N552, N588);
nor NOR2_229 (N661, N587, N589);
not NOT1_230 (N662, N590);
and AND2_231 (N665, N593, N590);
nor NOR2_232 (N669, N596, N522);
not NOT1_233 (N670, N597);
and AND2_234 (N673, N600, N597);
nor NOR2_235 (N677, N605, N523);
not NOT1_236 (N678, N606);
and AND2_237 (N682, N609, N606);
nor NOR2_238 (N686, N615, N524);
not NOT1_239 (N687, N616);
and AND2_240 (N692, N619, N616);
nor NOR2_241 (N696, N624, N525);
not NOT1_242 (N697, N625);
and AND2_243 (N700, N628, N625);
nor NOR2_244 (N704, N631, N526);
not NOT1_245 (N705, N632);
and AND2_246 (N708, N635, N632);
nor NOR2_247 (N712, N337, N640);
not NOT1_248 (N713, N641);
and AND2_249 (N717, N644, N641);
nor NOR2_250 (N721, N339, N650);
not NOT1_251 (N722, N651);
and AND2_252 (N727, N654, N651);
nor NOR2_253 (N731, N341, N659);
nand NAND2_254 (N732, N654, N261);
nand NAND3_255 (N733, N644, N654, N261);
nand NAND4_256 (N734, N635, N644, N654, N261);
not NOT1_257 (N735, N662);
and AND2_258 (N736, N228, N665);
and AND2_259 (N737, N237, N662);
not NOT1_260 (N738, N670);
and AND2_261 (N739, N228, N673);
and AND2_262 (N740, N237, N670);
not NOT1_263 (N741, N678);
and AND2_264 (N742, N228, N682);
and AND2_265 (N743, N237, N678);
not NOT1_266 (N744, N687);
and AND2_267 (N745, N228, N692);
and AND2_268 (N746, N237, N687);
not NOT1_269 (N747, N697);
and AND2_270 (N748, N228, N700);
and AND2_271 (N749, N237, N697);
not NOT1_272 (N750, N705);
and AND2_273 (N751, N228, N708);
and AND2_274 (N752, N237, N705);
not NOT1_275 (N753, N713);
and AND2_276 (N754, N228, N717);
and AND2_277 (N755, N237, N713);
not NOT1_278 (N756, N722);
nor NOR2_279 (N757, N727, N261);
and AND2_280 (N758, N727, N261);
and AND2_281 (N759, N228, N727);
and AND2_282 (N760, N237, N722);
nand NAND2_283 (N761, N644, N722);
nand NAND2_284 (N762, N635, N713);
nand NAND3_285 (N763, N635, N644, N722);
nand NAND2_286 (N764, N609, N687);
nand NAND2_287 (N765, N600, N678);
nand NAND3_288 (N766, N600, N609, N687);
buf BUFF1_289 (N767, N660);
buf BUFF1_290 (N768, N661);
nor NOR2_291 (N769, N736, N737);
nor NOR2_292 (N770, N739, N740);
nor NOR2_293 (N771, N742, N743);
nor NOR2_294 (N772, N745, N746);
nand NAND4_295 (N773, N750, N762, N763, N734);
nor NOR2_296 (N777, N748, N749);
nand NAND3_297 (N778, N753, N761, N733);
nor NOR2_298 (N781, N751, N752);
nand NAND2_299 (N782, N756, N732);
nor NOR2_300 (N785, N754, N755);
nor NOR2_301 (N786, N757, N758);
nor NOR2_302 (N787, N759, N760);
nor NOR2_303 (N788, N700, N773);
and AND2_304 (N789, N700, N773);
nor NOR2_305 (N790, N708, N778);
and AND2_306 (N791, N708, N778);
nor NOR2_307 (N792, N717, N782);
and AND2_308 (N793, N717, N782);
and AND2_309 (N794, N219, N786);
nand NAND2_310 (N795, N628, N773);
nand NAND2_311 (N796, N795, N747);
nor NOR2_312 (N802, N788, N789);
nor NOR2_313 (N803, N790, N791);
nor NOR2_314 (N804, N792, N793);
nor NOR2_315 (N805, N340, N794);
nor NOR2_316 (N806, N692, N796);
and AND2_317 (N807, N692, N796);
and AND2_318 (N808, N219, N802);
and AND2_319 (N809, N219, N803);
and AND2_320 (N810, N219, N804);
nand NAND4_321 (N811, N805, N787, N731, N529);
nand NAND2_322 (N812, N619, N796);
nand NAND3_323 (N813, N609, N619, N796);
nand NAND4_324 (N814, N600, N609, N619, N796);
nand NAND4_325 (N815, N738, N765, N766, N814);
nand NAND3_326 (N819, N741, N764, N813);
nand NAND2_327 (N822, N744, N812);
nor NOR2_328 (N825, N806, N807);
nor NOR2_329 (N826, N335, N808);
nor NOR2_330 (N827, N336, N809);
nor NOR2_331 (N828, N338, N810);
not NOT1_332 (N829, N811);
nor NOR2_333 (N830, N665, N815);
and AND2_334 (N831, N665, N815);
nor NOR2_335 (N832, N673, N819);
and AND2_336 (N833, N673, N819);
nor NOR2_337 (N834, N682, N822);
and AND2_338 (N835, N682, N822);
and AND2_339 (N836, N219, N825);
nand NAND3_340 (N837, N826, N777, N704);
nand NAND4_341 (N838, N827, N781, N712, N527);
nand NAND4_342 (N839, N828, N785, N721, N528);
not NOT1_343 (N840, N829);
nand NAND2_344 (N841, N815, N593);
nor NOR2_345 (N842, N830, N831);
nor NOR2_346 (N843, N832, N833);
nor NOR2_347 (N844, N834, N835);
nor NOR2_348 (N845, N334, N836);
not NOT1_349 (N846, N837);
not NOT1_350 (N847, N838);
not NOT1_351 (N848, N839);
and AND2_352 (N849, N735, N841);
buf BUFF1_353 (N850, N840);
and AND2_354 (N851, N219, N842);
and AND2_355 (N852, N219, N843);
and AND2_356 (N853, N219, N844);
nand NAND3_357 (N854, N845, N772, N696);
not NOT1_358 (N855, N846);
not NOT1_359 (N856, N847);
not NOT1_360 (N857, N848);
not NOT1_361 (N858, N849);
nor NOR2_362 (N859, N417, N851);
nor NOR2_363 (N860, N332, N852);
nor NOR2_364 (N861, N333, N853);
not NOT1_365 (N862, N854);
buf BUFF1_366 (N863, N855);
buf BUFF1_367 (N864, N856);
buf BUFF1_368 (N865, N857);
buf BUFF1_369 (N866, N858);
nand NAND3_370 (N867, N859, N769, N669);
nand NAND3_371 (N868, N860, N770, N677);
nand NAND3_372 (N869, N861, N771, N686);
not NOT1_373 (N870, N862);
not NOT1_374 (N871, N867);
not NOT1_375 (N872, N868);
not NOT1_376 (N873, N869);
buf BUFF1_377 (N874, N870);
not NOT1_378 (N875, N871);
not NOT1_379 (N876, N872);
not NOT1_380 (N877, N873);
buf BUFF1_381 (N878, N875);
buf BUFF1_382 (N879, N876);
buf BUFF1_383 (N880, N877);

endmodule




//OUTPUT

/*(base) bhaavanaa@bhaavanaa:~/VLSI_lab/DA2$ python da2.py 
enter the verilog file name: c880a.v

number of inputs=  60
inputs are:  ['N1', 'N8', 'N13', 'N17', 'N26', 'N29', 'N36', 'N42', 'N51', 'N55', 'N59', 'N68', 'N72', 'N73', 'N74', 'N75', 'N80', 'N85', 'N86', 'N87', 'N88', 'N89', 'N90', 'N91', 'N96', 'N101', 'N106', 'N111', 'N116', 'N121', 'N126', 'N130', 'N135', 'N138', 'N143', 'N146', 'N149', 'N152', 'N153', 'N156', 'N159', 'N165', 'N171', 'N177', 'N183', 'N189', 'N195', 'N201', 'N207', 'N210', 'N219', 'N228', 'N237', 'N246', 'N255', 'N259', 'N260', 'N261', 'N267', 'N268']



number of wires=  357
intermediate wires are:  ['N269', 'N270', 'N273', 'N276', 'N279', 'N280', 'N284', 'N285', 'N286', 'N287', 'N290', 'N291', 'N292', 'N293', 'N294', 'N295', 'N296', 'N297', 'N298', 'N301', 'N302', 'N303', 'N304', 'N305', 'N306', 'N307', 'N308', 'N309', 'N310', 'N316', 'N317', 'N318', 'N319', 'N322', 'N323', 'N324', 'N325', 'N326', 'N327', 'N328', 'N329', 'N330', 'N331', 'N332', 'N333', 'N334', 'N335', 'N336', 'N337', 'N338', 'N339', 'N340', 'N341', 'N342', 'N343', 'N344', 'N345', 'N346', 'N347', 'N348', 'N349', 'N350', 'N351', 'N352', 'N353', 'N354', 'N355', 'N356', 'N357', 'N360', 'N363', 'N366', 'N369', 'N375', 'N376', 'N379', 'N382', 'N385', 'N392', 'N393', 'N399', 'N400', 'N401', 'N402', 'N403', 'N404', 'N405', 'N406', 'N407', 'N408', 'N409', 'N410', 'N411', 'N412', 'N413', 'N414', 'N415', 'N416', 'N417', 'N424', 'N425', 'N426', 'N427', 'N432', 'N437', 'N442', 'N443', 'N444', 'N445', 'N451', 'N460', 'N463', 'N466', 'N475', 'N476', 'N477', 'N478', 'N479', 'N480', 'N481', 'N482', 'N483', 'N488', 'N489', 'N490', 'N491', 'N492', 'N495', 'N498', 'N499', 'N500', 'N501', 'N502', 'N503', 'N504', 'N505', 'N506', 'N507', 'N508', 'N509', 'N510', 'N511', 'N512', 'N513', 'N514', 'N515', 'N516', 'N517', 'N518', 'N519', 'N520', 'N521', 'N522', 'N523', 'N524', 'N525', 'N526', 'N527', 'N528', 'N529', 'N530', 'N533', 'N536', 'N537', 'N538', 'N539', 'N540', 'N541', 'N542', 'N543', 'N544', 'N547', 'N550', 'N551', 'N552', 'N553', 'N557', 'N561', 'N565', 'N569', 'N573', 'N577', 'N581', 'N585', 'N586', 'N587', 'N588', 'N589', 'N590', 'N593', 'N596', 'N597', 'N600', 'N605', 'N606', 'N609', 'N615', 'N616', 'N619', 'N624', 'N625', 'N628', 'N631', 'N632', 'N635', 'N640', 'N641', 'N644', 'N650', 'N651', 'N654', 'N659', 'N660', 'N661', 'N662', 'N665', 'N669', 'N670', 'N673', 'N677', 'N678', 'N682', 'N686', 'N687', 'N692', 'N696', 'N697', 'N700', 'N704', 'N705', 'N708', 'N712', 'N713', 'N717', 'N721', 'N722', 'N727', 'N731', 'N732', 'N733', 'N734', 'N735', 'N736', 'N737', 'N738', 'N739', 'N740', 'N741', 'N742', 'N743', 'N744', 'N745', 'N746', 'N747', 'N748', 'N749', 'N750', 'N751', 'N752', 'N753', 'N754', 'N755', 'N756', 'N757', 'N758', 'N759', 'N760', 'N761', 'N762', 'N763', 'N764', 'N765', 'N766', 'N769', 'N770', 'N771', 'N772', 'N773', 'N777', 'N778', 'N781', 'N782', 'N785', 'N786', 'N787', 'N788', 'N789', 'N790', 'N791', 'N792', 'N793', 'N794', 'N795', 'N796', 'N802', 'N803', 'N804', 'N805', 'N806', 'N807', 'N808', 'N809', 'N810', 'N811', 'N812', 'N813', 'N814', 'N815', 'N819', 'N822', 'N825', 'N826', 'N827', 'N828', 'N829', 'N830', 'N831', 'N832', 'N833', 'N834', 'N835', 'N836', 'N837', 'N838', 'N839', 'N840', 'N841', 'N842', 'N843', 'N844', 'N845', 'N846', 'N847', 'N848', 'N849', 'N851', 'N852', 'N853', 'N854', 'N855', 'N856', 'N857', 'N858', 'N859', 'N860', 'N861', 'N862', 'N867', 'N868', 'N869', 'N870', 'N871', 'N872', 'N873', 'N875', 'N876', 'N877']



number of outputs=  26
outputs are:  ['N388', 'N389', 'N390', 'N391', 'N418', 'N419', 'N420', 'N421', 'N422', 'N423', 'N446', 'N447', 'N448', 'N449', 'N450', 'N767', 'N768', 'N850', 'N863', 'N864', 'N865', 'N866', 'N874', 'N878', 'N879', 'N880']



number of gates=  383
gate array is:  [['nand', 'N269', 'N1', 'N8', 'N13', 'N17'], ['nand', 'N270', 'N1', 'N26', 'N13', 'N17'], ['and', 'N273', 'N29', 'N36', 'N42'], ['and', 'N276', 'N1', 'N26', 'N51'], ['nand', 'N279', 'N1', 'N8', 'N51', 'N17'], ['nand', 'N280', 'N1', 'N8', 'N13', 'N55'], ['nand', 'N284', 'N59', 'N42', 'N68', 'N72'], ['nand', 'N285', 'N29', 'N68'], ['nand', 'N286', 'N59', 'N68', 'N74'], ['and', 'N287', 'N29', 'N75', 'N80'], ['and', 'N290', 'N29', 'N75', 'N42'], ['and', 'N291', 'N29', 'N36', 'N80'], ['and', 'N292', 'N29', 'N36', 'N42'], ['and', 'N293', 'N59', 'N75', 'N80'], ['and', 'N294', 'N59', 'N75', 'N42'], ['and', 'N295', 'N59', 'N36', 'N80'], ['and', 'N296', 'N59', 'N36', 'N42'], ['and', 'N297', 'N85', 'N86'], ['or', 'N298', 'N87', 'N88'], ['nand', 'N301', 'N91', 'N96'], ['or', 'N302', 'N91', 'N96'], ['nand', 'N303', 'N101', 'N106'], ['or', 'N304', 'N101', 'N106'], ['nand', 'N305', 'N111', 'N116'], ['or', 'N306', 'N111', 'N116'], ['nand', 'N307', 'N121', 'N126'], ['or', 'N308', 'N121', 'N126'], ['and', 'N309', 'N8', 'N138'], ['not', 'N310', 'N268'], ['and', 'N316', 'N51', 'N138'], ['and', 'N317', 'N17', 'N138'], ['and', 'N318', 'N152', 'N138'], ['nand', 'N319', 'N59', 'N156'], ['nor', 'N322', 'N17', 'N42'], ['and', 'N323', 'N17', 'N42'], ['nand', 'N324', 'N159', 'N165'], ['or', 'N325', 'N159', 'N165'], ['nand', 'N326', 'N171', 'N177'], ['or', 'N327', 'N171', 'N177'], ['nand', 'N328', 'N183', 'N189'], ['or', 'N329', 'N183', 'N189'], ['nand', 'N330', 'N195', 'N201'], ['or', 'N331', 'N195', 'N201'], ['and', 'N332', 'N210', 'N91'], ['and', 'N333', 'N210', 'N96'], ['and', 'N334', 'N210', 'N101'], ['and', 'N335', 'N210', 'N106'], ['and', 'N336', 'N210', 'N111'], ['and', 'N337', 'N255', 'N259'], ['and', 'N338', 'N210', 'N116'], ['and', 'N339', 'N255', 'N260'], ['and', 'N340', 'N210', 'N121'], ['and', 'N341', 'N255', 'N267'], ['not', 'N342', 'N269'], ['not', 'N343', 'N273'], ['or', 'N344', 'N270', 'N273'], ['not', 'N345', 'N276'], ['not', 'N346', 'N276'], ['not', 'N347', 'N279'], ['nor', 'N348', 'N280', 'N284'], ['or', 'N349', 'N280', 'N285'], ['or', 'N350', 'N280', 'N286'], ['not', 'N351', 'N293'], ['not', 'N352', 'N294'], ['not', 'N353', 'N295'], ['not', 'N354', 'N296'], ['nand', 'N355', 'N89', 'N298'], ['and', 'N356', 'N90', 'N298'], ['nand', 'N357', 'N301', 'N302'], ['nand', 'N360', 'N303', 'N304'], ['nand', 'N363', 'N305', 'N306'], ['nand', 'N366', 'N307', 'N308'], ['not', 'N369', 'N310'], ['nor', 'N375', 'N322', 'N323'], ['nand', 'N376', 'N324', 'N325'], ['nand', 'N379', 'N326', 'N327'], ['nand', 'N382', 'N328', 'N329'], ['nand', 'N385', 'N330', 'N331'], ['buf', 'N388', 'N290'], ['buf', 'N389', 'N291'], ['buf', 'N390', 'N292'], ['buf', 'N391', 'N297'], ['or', 'N392', 'N270', 'N343'], ['not', 'N393', 'N345'], ['not', 'N399', 'N346'], ['and', 'N400', 'N348', 'N73'], ['not', 'N401', 'N349'], ['not', 'N402', 'N350'], ['not', 'N403', 'N355'], ['not', 'N404', 'N357'], ['not', 'N405', 'N360'], ['and', 'N406', 'N357', 'N360'], ['not', 'N407', 'N363'], ['not', 'N408', 'N366'], ['and', 'N409', 'N363', 'N366'], ['nand', 'N410', 'N347', 'N352'], ['not', 'N411', 'N376'], ['not', 'N412', 'N379'], ['and', 'N413', 'N376', 'N379'], ['not', 'N414', 'N382'], ['not', 'N415', 'N385'], ['and', 'N416', 'N382', 'N385'], ['and', 'N417', 'N210', 'N369'], ['buf', 'N418', 'N342'], ['buf', 'N419', 'N344'], ['buf', 'N420', 'N351'], ['buf', 'N421', 'N353'], ['buf', 'N422', 'N354'], ['buf', 'N423', 'N356'], ['not', 'N424', 'N400'], ['and', 'N425', 'N404', 'N405'], ['and', 'N426', 'N407', 'N408'], ['and', 'N427', 'N319', 'N393', 'N55'], ['and', 'N432', 'N393', 'N17', 'N287'], ['nand', 'N437', 'N393', 'N287', 'N55'], ['nand', 'N442', 'N375', 'N59', 'N156', 'N393'], ['nand', 'N443', 'N393', 'N319', 'N17'], ['and', 'N444', 'N411', 'N412'], ['and', 'N445', 'N414', 'N415'], ['buf', 'N446', 'N392'], ['buf', 'N447', 'N399'], ['buf', 'N448', 'N401'], ['buf', 'N449', 'N402'], ['buf', 'N450', 'N403'], ['not', 'N451', 'N424'], ['nor', 'N460', 'N406', 'N425'], ['nor', 'N463', 'N409', 'N426'], ['nand', 'N466', 'N442', 'N410'], ['and', 'N475', 'N143', 'N427'], ['and', 'N476', 'N310', 'N432'], ['and', 'N477', 'N146', 'N427'], ['and', 'N478', 'N310', 'N432'], ['and', 'N479', 'N149', 'N427'], ['and', 'N480', 'N310', 'N432'], ['and', 'N481', 'N153', 'N427'], ['and', 'N482', 'N310', 'N432'], ['nand', 'N483', 'N443', 'N1'], ['or', 'N488', 'N369', 'N437'], ['or', 'N489', 'N369', 'N437'], ['or', 'N490', 'N369', 'N437'], ['or', 'N491', 'N369', 'N437'], ['nor', 'N492', 'N413', 'N444'], ['nor', 'N495', 'N416', 'N445'], ['nand', 'N498', 'N130', 'N460'], ['or', 'N499', 'N130', 'N460'], ['nand', 'N500', 'N463', 'N135'], ['or', 'N501', 'N463', 'N135'], ['and', 'N502', 'N91', 'N466'], ['nor', 'N503', 'N475', 'N476'], ['and', 'N504', 'N96', 'N466'], ['nor', 'N505', 'N477', 'N478'], ['and', 'N506', 'N101', 'N466'], ['nor', 'N507', 'N479', 'N480'], ['and', 'N508', 'N106', 'N466'], ['nor', 'N509', 'N481', 'N482'], ['and', 'N510', 'N143', 'N483'], ['and', 'N511', 'N111', 'N466'], ['and', 'N512', 'N146', 'N483'], ['and', 'N513', 'N116', 'N466'], ['and', 'N514', 'N149', 'N483'], ['and', 'N515', 'N121', 'N466'], ['and', 'N516', 'N153', 'N483'], ['and', 'N517', 'N126', 'N466'], ['nand', 'N518', 'N130', 'N492'], ['or', 'N519', 'N130', 'N492'], ['nand', 'N520', 'N495', 'N207'], ['or', 'N521', 'N495', 'N207'], ['and', 'N522', 'N451', 'N159'], ['and', 'N523', 'N451', 'N165'], ['and', 'N524', 'N451', 'N171'], ['and', 'N525', 'N451', 'N177'], ['and', 'N526', 'N451', 'N183'], ['nand', 'N527', 'N451', 'N189'], ['nand', 'N528', 'N451', 'N195'], ['nand', 'N529', 'N451', 'N201'], ['nand', 'N530', 'N498', 'N499'], ['nand', 'N533', 'N500', 'N501'], ['nor', 'N536', 'N309', 'N502'], ['nor', 'N537', 'N316', 'N504'], ['nor', 'N538', 'N317', 'N506'], ['nor', 'N539', 'N318', 'N508'], ['nor', 'N540', 'N510', 'N511'], ['nor', 'N541', 'N512', 'N513'], ['nor', 'N542', 'N514', 'N515'], ['nor', 'N543', 'N516', 'N517'], ['nand', 'N544', 'N518', 'N519'], ['nand', 'N547', 'N520', 'N521'], ['not', 'N550', 'N530'], ['not', 'N551', 'N533'], ['and', 'N552', 'N530', 'N533'], ['nand', 'N553', 'N536', 'N503'], ['nand', 'N557', 'N537', 'N505'], ['nand', 'N561', 'N538', 'N507'], ['nand', 'N565', 'N539', 'N509'], ['nand', 'N569', 'N488', 'N540'], ['nand', 'N573', 'N489', 'N541'], ['nand', 'N577', 'N490', 'N542'], ['nand', 'N581', 'N491', 'N543'], ['not', 'N585', 'N544'], ['not', 'N586', 'N547'], ['and', 'N587', 'N544', 'N547'], ['and', 'N588', 'N550', 'N551'], ['and', 'N589', 'N585', 'N586'], ['nand', 'N590', 'N553', 'N159'], ['or', 'N593', 'N553', 'N159'], ['and', 'N596', 'N246', 'N553'], ['nand', 'N597', 'N557', 'N165'], ['or', 'N600', 'N557', 'N165'], ['and', 'N605', 'N246', 'N557'], ['nand', 'N606', 'N561', 'N171'], ['or', 'N609', 'N561', 'N171'], ['and', 'N615', 'N246', 'N561'], ['nand', 'N616', 'N565', 'N177'], ['or', 'N619', 'N565', 'N177'], ['and', 'N624', 'N246', 'N565'], ['nand', 'N625', 'N569', 'N183'], ['or', 'N628', 'N569', 'N183'], ['and', 'N631', 'N246', 'N569'], ['nand', 'N632', 'N573', 'N189'], ['or', 'N635', 'N573', 'N189'], ['and', 'N640', 'N246', 'N573'], ['nand', 'N641', 'N577', 'N195'], ['or', 'N644', 'N577', 'N195'], ['and', 'N650', 'N246', 'N577'], ['nand', 'N651', 'N581', 'N201'], ['or', 'N654', 'N581', 'N201'], ['and', 'N659', 'N246', 'N581'], ['nor', 'N660', 'N552', 'N588'], ['nor', 'N661', 'N587', 'N589'], ['not', 'N662', 'N590'], ['and', 'N665', 'N593', 'N590'], ['nor', 'N669', 'N596', 'N522'], ['not', 'N670', 'N597'], ['and', 'N673', 'N600', 'N597'], ['nor', 'N677', 'N605', 'N523'], ['not', 'N678', 'N606'], ['and', 'N682', 'N609', 'N606'], ['nor', 'N686', 'N615', 'N524'], ['not', 'N687', 'N616'], ['and', 'N692', 'N619', 'N616'], ['nor', 'N696', 'N624', 'N525'], ['not', 'N697', 'N625'], ['and', 'N700', 'N628', 'N625'], ['nor', 'N704', 'N631', 'N526'], ['not', 'N705', 'N632'], ['and', 'N708', 'N635', 'N632'], ['nor', 'N712', 'N337', 'N640'], ['not', 'N713', 'N641'], ['and', 'N717', 'N644', 'N641'], ['nor', 'N721', 'N339', 'N650'], ['not', 'N722', 'N651'], ['and', 'N727', 'N654', 'N651'], ['nor', 'N731', 'N341', 'N659'], ['nand', 'N732', 'N654', 'N261'], ['nand', 'N733', 'N644', 'N654', 'N261'], ['nand', 'N734', 'N635', 'N644', 'N654', 'N261'], ['not', 'N735', 'N662'], ['and', 'N736', 'N228', 'N665'], ['and', 'N737', 'N237', 'N662'], ['not', 'N738', 'N670'], ['and', 'N739', 'N228', 'N673'], ['and', 'N740', 'N237', 'N670'], ['not', 'N741', 'N678'], ['and', 'N742', 'N228', 'N682'], ['and', 'N743', 'N237', 'N678'], ['not', 'N744', 'N687'], ['and', 'N745', 'N228', 'N692'], ['and', 'N746', 'N237', 'N687'], ['not', 'N747', 'N697'], ['and', 'N748', 'N228', 'N700'], ['and', 'N749', 'N237', 'N697'], ['not', 'N750', 'N705'], ['and', 'N751', 'N228', 'N708'], ['and', 'N752', 'N237', 'N705'], ['not', 'N753', 'N713'], ['and', 'N754', 'N228', 'N717'], ['and', 'N755', 'N237', 'N713'], ['not', 'N756', 'N722'], ['nor', 'N757', 'N727', 'N261'], ['and', 'N758', 'N727', 'N261'], ['and', 'N759', 'N228', 'N727'], ['and', 'N760', 'N237', 'N722'], ['nand', 'N761', 'N644', 'N722'], ['nand', 'N762', 'N635', 'N713'], ['nand', 'N763', 'N635', 'N644', 'N722'], ['nand', 'N764', 'N609', 'N687'], ['nand', 'N765', 'N600', 'N678'], ['nand', 'N766', 'N600', 'N609', 'N687'], ['buf', 'N767', 'N660'], ['buf', 'N768', 'N661'], ['nor', 'N769', 'N736', 'N737'], ['nor', 'N770', 'N739', 'N740'], ['nor', 'N771', 'N742', 'N743'], ['nor', 'N772', 'N745', 'N746'], ['nand', 'N773', 'N750', 'N762', 'N763', 'N734'], ['nor', 'N777', 'N748', 'N749'], ['nand', 'N778', 'N753', 'N761', 'N733'], ['nor', 'N781', 'N751', 'N752'], ['nand', 'N782', 'N756', 'N732'], ['nor', 'N785', 'N754', 'N755'], ['nor', 'N786', 'N757', 'N758'], ['nor', 'N787', 'N759', 'N760'], ['nor', 'N788', 'N700', 'N773'], ['and', 'N789', 'N700', 'N773'], ['nor', 'N790', 'N708', 'N778'], ['and', 'N791', 'N708', 'N778'], ['nor', 'N792', 'N717', 'N782'], ['and', 'N793', 'N717', 'N782'], ['and', 'N794', 'N219', 'N786'], ['nand', 'N795', 'N628', 'N773'], ['nand', 'N796', 'N795', 'N747'], ['nor', 'N802', 'N788', 'N789'], ['nor', 'N803', 'N790', 'N791'], ['nor', 'N804', 'N792', 'N793'], ['nor', 'N805', 'N340', 'N794'], ['nor', 'N806', 'N692', 'N796'], ['and', 'N807', 'N692', 'N796'], ['and', 'N808', 'N219', 'N802'], ['and', 'N809', 'N219', 'N803'], ['and', 'N810', 'N219', 'N804'], ['nand', 'N811', 'N805', 'N787', 'N731', 'N529'], ['nand', 'N812', 'N619', 'N796'], ['nand', 'N813', 'N609', 'N619', 'N796'], ['nand', 'N814', 'N600', 'N609', 'N619', 'N796'], ['nand', 'N815', 'N738', 'N765', 'N766', 'N814'], ['nand', 'N819', 'N741', 'N764', 'N813'], ['nand', 'N822', 'N744', 'N812'], ['nor', 'N825', 'N806', 'N807'], ['nor', 'N826', 'N335', 'N808'], ['nor', 'N827', 'N336', 'N809'], ['nor', 'N828', 'N338', 'N810'], ['not', 'N829', 'N811'], ['nor', 'N830', 'N665', 'N815'], ['and', 'N831', 'N665', 'N815'], ['nor', 'N832', 'N673', 'N819'], ['and', 'N833', 'N673', 'N819'], ['nor', 'N834', 'N682', 'N822'], ['and', 'N835', 'N682', 'N822'], ['and', 'N836', 'N219', 'N825'], ['nand', 'N837', 'N826', 'N777', 'N704'], ['nand', 'N838', 'N827', 'N781', 'N712', 'N527'], ['nand', 'N839', 'N828', 'N785', 'N721', 'N528'], ['not', 'N840', 'N829'], ['nand', 'N841', 'N815', 'N593'], ['nor', 'N842', 'N830', 'N831'], ['nor', 'N843', 'N832', 'N833'], ['nor', 'N844', 'N834', 'N835'], ['nor', 'N845', 'N334', 'N836'], ['not', 'N846', 'N837'], ['not', 'N847', 'N838'], ['not', 'N848', 'N839'], ['and', 'N849', 'N735', 'N841'], ['buf', 'N850', 'N840'], ['and', 'N851', 'N219', 'N842'], ['and', 'N852', 'N219', 'N843'], ['and', 'N853', 'N219', 'N844'], ['nand', 'N854', 'N845', 'N772', 'N696'], ['not', 'N855', 'N846'], ['not', 'N856', 'N847'], ['not', 'N857', 'N848'], ['not', 'N858', 'N849'], ['nor', 'N859', 'N417', 'N851'], ['nor', 'N860', 'N332', 'N852'], ['nor', 'N861', 'N333', 'N853'], ['not', 'N862', 'N854'], ['buf', 'N863', 'N855'], ['buf', 'N864', 'N856'], ['buf', 'N865', 'N857'], ['buf', 'N866', 'N858'], ['nand', 'N867', 'N859', 'N769', 'N669'], ['nand', 'N868', 'N860', 'N770', 'N677'], ['nand', 'N869', 'N861', 'N771', 'N686'], ['not', 'N870', 'N862'], ['not', 'N871', 'N867'], ['not', 'N872', 'N868'], ['not', 'N873', 'N869'], ['buf', 'N874', 'N870'], ['not', 'N875', 'N871'], ['not', 'N876', 'N872'], ['not', 'N877', 'N873'], ['buf', 'N878', 'N875'], ['buf', 'N879', 'N876'], ['buf', 'N880', 'N877']]


input probabilities: 
N1 0.5
N8 0.5
N13 0.5
N17 0.5
N26 0.5
N29 0.5
N36 0.5
N42 0.5
N51 0.5
N55 0.5
N59 0.5
N68 0.5
N72 0.5
N73 0.5
N74 0.5
N75 0.5
N80 0.5
N85 0.5
N86 0.5
N87 0.5
N88 0.5
N89 0.5
N90 0.5
N91 0.5
N96 0.5
N101 0.5
N106 0.5
N111 0.5
N116 0.5
N121 0.5
N126 0.5
N130 0.5
N135 0.5
N138 0.5
N143 0.5
N146 0.5
N149 0.5
N152 0.5
N153 0.5
N156 0.5
N159 0.5
N165 0.5
N171 0.5
N177 0.5
N183 0.5
N189 0.5
N195 0.5
N201 0.5
N207 0.5
N210 0.5
N219 0.5
N228 0.5
N237 0.5
N246 0.5
N255 0.5
N259 0.5
N260 0.5
N261 0.5
N267 0.5
N268 0.5


probability of intermediate wires:
N269 0.9375
N270 0.9375
N273 0.125
N276 0.125
N279 0.9375
N280 0.9375
N284 0.9375
N285 0.75
N286 0.875
N287 0.125
N290 0.125
N291 0.125
N292 0.125
N293 0.125
N294 0.125
N295 0.125
N296 0.125
N297 0.25
N298 0.75
N301 0.75
N302 0.75
N303 0.75
N304 0.75
N305 0.75
N306 0.75
N307 0.75
N308 0.75
N309 0.25
N310 0.5
N316 0.25
N317 0.25
N318 0.25
N319 0.75
N322 0.25
N323 0.25
N324 0.75
N325 0.75
N326 0.75
N327 0.75
N328 0.75
N329 0.75
N330 0.75
N331 0.75
N332 0.25
N333 0.25
N334 0.25
N335 0.25
N336 0.25
N337 0.25
N338 0.25
N339 0.25
N340 0.25
N341 0.25
N342 0.0625
N343 0.875
N344 0.9453125
N345 0.875
N346 0.875
N347 0.0625
N348 0.00390625
N349 0.984375
N350 0.9921875
N351 0.875
N352 0.875
N353 0.875
N354 0.875
N355 0.625
N356 0.375
N357 0.4375
N360 0.4375
N363 0.4375
N366 0.4375
N369 0.5
N375 0.5625
N376 0.4375
N379 0.4375
N382 0.4375
N385 0.4375
N392 0.9921875
N393 0.125
N399 0.125
N400 0.001953125
N401 0.015625
N402 0.0078125
N403 0.375
N404 0.5625
N405 0.5625
N406 0.19140625
N407 0.5625
N408 0.5625
N409 0.19140625
N410 0.9453125
N411 0.5625
N412 0.5625
N413 0.19140625
N414 0.5625
N415 0.5625
N416 0.19140625
N417 0.25
N424 0.998046875
N425 0.31640625
N426 0.31640625
N427 0.046875
N432 0.0078125
N437 0.9921875
N442 0.982421875
N443 0.953125
N444 0.31640625
N445 0.31640625
N451 0.001953125
N460 0.5527496337890625
N463 0.5527496337890625
N466 0.0713043212890625
N475 0.0234375
N476 0.00390625
N477 0.0234375
N478 0.00390625
N479 0.0234375
N480 0.00390625
N481 0.0234375
N482 0.00390625
N483 0.5234375
N488 0.99609375
N489 0.99609375
N490 0.99609375
N491 0.99609375
N492 0.5527496337890625
N495 0.5527496337890625
N498 0.7236251831054688
N499 0.7763748168945312
N500 0.7236251831054688
N501 0.7763748168945312
N502 0.03565216064453125
N503 0.972747802734375
N504 0.03565216064453125
N505 0.972747802734375
N506 0.03565216064453125
N507 0.972747802734375
N508 0.03565216064453125
N509 0.972747802734375
N510 0.26171875
N511 0.03565216064453125
N512 0.26171875
N513 0.03565216064453125
N514 0.26171875
N515 0.03565216064453125
N516 0.26171875
N517 0.03565216064453125
N518 0.7236251831054688
N519 0.7763748168945312
N520 0.7236251831054688
N521 0.7763748168945312
N522 0.0009765625
N523 0.0009765625
N524 0.0009765625
N525 0.0009765625
N526 0.0009765625
N527 0.9990234375
N528 0.9990234375
N529 0.9990234375
N530 0.43819563096622005
N533 0.43819563096622005
N536 0.7232608795166016
N537 0.7232608795166016
N538 0.7232608795166016
N539 0.7232608795166016
N540 0.7119599282741547
N541 0.7119599282741547
N542 0.7119599282741547
N543 0.7119599282741547
N544 0.43819563096622005
N547 0.43819563096622005
N550 0.56180436903378
N551 0.56180436903378
N552 0.19201541099788372
N553 0.2964495686464943
N557 0.2964495686464943
N561 0.2964495686464943
N565 0.2964495686464943
N569 0.29082116519566625
N573 0.29082116519566625
N577 0.29082116519566625
N581 0.29082116519566625
N585 0.56180436903378
N586 0.56180436903378
N587 0.19201541099788372
N588 0.3156241490654436
N589 0.3156241490654436
N590 0.8517752156767529
N593 0.6482247843232471
N596 0.14822478432324715
N597 0.8517752156767529
N600 0.6482247843232471
N605 0.14822478432324715
N606 0.8517752156767529
N609 0.6482247843232471
N615 0.14822478432324715
N616 0.8517752156767529
N619 0.6482247843232471
N624 0.14822478432324715
N625 0.8545894174021669
N628 0.6454105825978331
N631 0.14541058259783313
N632 0.8545894174021669
N635 0.6454105825978331
N640 0.14541058259783313
N641 0.8545894174021669
N644 0.6454105825978331
N650 0.14541058259783313
N651 0.8545894174021669
N654 0.6454105825978331
N659 0.14541058259783313
N660 0.5529651406403311
N661 0.5529651406403311
N662 0.14822478432324715
N665 0.5521418054739504
N669 0.8509434039426935
N670 0.14822478432324715
N673 0.5521418054739504
N677 0.8509434039426935
N678 0.14822478432324715
N682 0.5521418054739504
N686 0.8509434039426935
N687 0.14822478432324715
N692 0.5521418054739504
N696 0.8509434039426935
N697 0.14541058259783313
N700 0.5515610537674753
N704 0.8537548574242351
N705 0.14541058259783313
N708 0.5515610537674753
N712 0.6409420630516252
N713 0.14541058259783313
N717 0.5515610537674753
N721 0.6409420630516252
N722 0.14541058259783313
N727 0.5515610537674753
N731 0.6409420630516252
N732 0.6772947087010834
N733 0.7917225899353628
N734 0.8655755554282147
N735 0.8517752156767529
N736 0.2760709027369752
N737 0.07411239216162357
N738 0.8517752156767529
N739 0.2760709027369752
N740 0.07411239216162357
N741 0.8517752156767529
N742 0.2760709027369752
N743 0.07411239216162357
N744 0.8517752156767529
N745 0.2760709027369752
N746 0.07411239216162357
N747 0.8545894174021669
N748 0.27578052688373766
N749 0.07270529129891656
N750 0.8545894174021669
N751 0.27578052688373766
N752 0.07270529129891656
N753 0.8545894174021669
N754 0.27578052688373766
N755 0.07270529129891656
N756 0.8545894174021669
N757 0.22421947311626234
N758 0.27578052688373766
N759 0.27578052688373766
N760 0.07270529129891656
N761 0.9061504711696422
N762 0.9061504711696422
N763 0.9394285209210667
N764 0.9039170211507033
N765 0.9039170211507033
N766 0.9377166317582795
N769 0.6702769801094574
N770 0.6702769801094574
N771 0.6702769801094574
N772 0.6702769801094574
N773 0.370310349418004
N777 0.6715648853589966
N778 0.38690063287509147
N781 0.6715648853589966
N782 0.4211911094815708
N785 0.6715648853589966
N786 0.5618353644335968
N787 0.6715648853589966
N788 0.28237736336051694
N789 0.20424876654599627
N790 0.27493763412932176
N791 0.21339932077188856
N792 0.25956044893410113
N793 0.23231261218314725
N794 0.2809176822167984
N795 0.7609977816401189
N796 0.34965934914382935
N802 0.5710490982603831
N803 0.570334549476617
N804 0.5684261047940631
N805 0.5393117383374011
N806 0.2912603897193406
N807 0.19306154433712033
N808 0.28552454913019154
N809 0.2851672747383085
N810 0.28421305239703154
N811 0.7680884899434697
N812 0.7733421438146343
N813 0.8530747600590717
N814 0.9047594180276504
N815 0.3467817722123865
N819 0.34318863903525043
N822 0.34128632866036746
N825 0.5719092465869865
N826 0.5358565881523564
N827 0.5361245439462686
N828 0.5368402107022263
N829 0.23191151005653032
N830 0.2925491361284664
N831 0.1914727138148033
N832 0.29415835026587017
N833 0.18948879477507102
N834 0.29501031555579343
N835 0.1884384496901113
N836 0.28595462329349325
N837 0.6927656697769178
N838 0.7694590276335446
N839 0.7691512810256493
N840 0.7680884899434697
N841 0.7752074605003924
N842 0.571993327075424
N843 0.5720925662239618
N844 0.5721425212600195
N845 0.5355340325298801
N846 0.3072343302230822
N847 0.23054097236645543
N848 0.23084871897435066
N849 0.6603025018619496
N851 0.285996663537712
N852 0.2860462831119809
N853 0.28607126063000976
N854 0.6945486454083917
N855 0.6927656697769178
N856 0.7694590276335446
N857 0.7691512810256493
N858 0.3396974981380504
N859 0.5355025023467159
N860 0.5354652876660143
N861 0.5354465545274927
N862 0.3054513545916083
N867 0.6945666292088095
N868 0.6945878552634401
N869 0.6945985400419781
N870 0.6945486454083917
N871 0.3054333707911905
N872 0.30541214473655987
N873 0.3054014599580219
N875 0.6945666292088095
N876 0.6945878552634401
N877 0.6945985400419781


probability of the outputs: 
N388 0.125
N389 0.125
N390 0.125
N391 0.25
N418 0.0625
N419 0.9453125
N420 0.875
N421 0.875
N422 0.875
N423 0.375
N446 0.9921875
N447 0.125
N448 0.015625
N449 0.0078125
N450 0.375
N767 0.5529651406403311
N768 0.5529651406403311
N850 0.7680884899434697
N863 0.6927656697769178
N864 0.7694590276335446
N865 0.7691512810256493
N866 0.3396974981380504
N874 0.6945486454083917
N878 0.6945666292088095
N879 0.6945878552634401
N880 0.6945985400419781


activity factors of intermediate wires:
N269 0.0586
N270 0.0586
N273 0.1094
N276 0.1094
N279 0.0586
N280 0.0586
N284 0.0586
N285 0.1875
N286 0.1094
N287 0.1094
N290 0.1094
N291 0.1094
N292 0.1094
N293 0.1094
N294 0.1094
N295 0.1094
N296 0.1094
N297 0.1875
N298 0.1875
N301 0.1875
N302 0.1875
N303 0.1875
N304 0.1875
N305 0.1875
N306 0.1875
N307 0.1875
N308 0.1875
N309 0.1875
N310 0.25
N316 0.1875
N317 0.1875
N318 0.1875
N319 0.1875
N322 0.1875
N323 0.1875
N324 0.1875
N325 0.1875
N326 0.1875
N327 0.1875
N328 0.1875
N329 0.1875
N330 0.1875
N331 0.1875
N332 0.1875
N333 0.1875
N334 0.1875
N335 0.1875
N336 0.1875
N337 0.1875
N338 0.1875
N339 0.1875
N340 0.1875
N341 0.1875
N342 0.0586
N343 0.1094
N344 0.0517
N345 0.1094
N346 0.1094
N347 0.0586
N348 0.0039
N349 0.0154
N350 0.0078
N351 0.1094
N352 0.1094
N353 0.1094
N354 0.1094
N355 0.2344
N356 0.2344
N357 0.2461
N360 0.2461
N363 0.2461
N366 0.2461
N369 0.25
N375 0.2461
N376 0.2461
N379 0.2461
N382 0.2461
N385 0.2461
N392 0.0078
N393 0.1094
N399 0.1094
N400 0.0019
N401 0.0154
N402 0.0078
N403 0.2344
N404 0.2461
N405 0.2461
N406 0.1548
N407 0.2461
N408 0.2461
N409 0.1548
N410 0.0517
N411 0.2461
N412 0.2461
N413 0.1548
N414 0.2461
N415 0.2461
N416 0.1548
N417 0.1875
N424 0.0019
N425 0.2163
N426 0.2163
N427 0.0447
N432 0.0078
N437 0.0078
N442 0.0173
N443 0.0447
N444 0.2163
N445 0.2163
N451 0.0019
N460 0.2472
N463 0.2472
N466 0.0662
N475 0.0229
N476 0.0039
N477 0.0229
N478 0.0039
N479 0.0229
N480 0.0039
N481 0.0229
N482 0.0039
N483 0.2495
N488 0.0039
N489 0.0039
N490 0.0039
N491 0.0039
N492 0.2472
N495 0.2472
N498 0.2
N499 0.1736
N500 0.2
N501 0.1736
N502 0.0344
N503 0.0265
N504 0.0344
N505 0.0265
N506 0.0344
N507 0.0265
N508 0.0344
N509 0.0265
N510 0.1932
N511 0.0344
N512 0.1932
N513 0.0344
N514 0.1932
N515 0.0344
N516 0.1932
N517 0.0344
N518 0.2
N519 0.1736
N520 0.2
N521 0.1736
N522 0.001
N523 0.001
N524 0.001
N525 0.001
N526 0.001
N527 0.001
N528 0.001
N529 0.001
N530 0.2462
N533 0.2462
N536 0.2002
N537 0.2002
N538 0.2002
N539 0.2002
N540 0.2051
N541 0.2051
N542 0.2051
N543 0.2051
N544 0.2462
N547 0.2462
N550 0.2462
N551 0.2462
N552 0.1551
N553 0.2086
N557 0.2086
N561 0.2086
N565 0.2086
N569 0.2062
N573 0.2062
N577 0.2062
N581 0.2062
N585 0.2462
N586 0.2462
N587 0.1551
N588 0.216
N589 0.216
N590 0.1263
N593 0.228
N596 0.1263
N597 0.1263
N600 0.228
N605 0.1263
N606 0.1263
N609 0.228
N615 0.1263
N616 0.1263
N619 0.228
N624 0.1263
N625 0.1243
N628 0.2289
N631 0.1243
N632 0.1243
N635 0.2289
N640 0.1243
N641 0.1243
N644 0.2289
N650 0.1243
N651 0.1243
N654 0.2289
N659 0.1243
N660 0.2472
N661 0.2472
N662 0.1263
N665 0.2473
N669 0.1268
N670 0.1263
N673 0.2473
N677 0.1268
N678 0.1263
N682 0.2473
N686 0.1268
N687 0.1263
N692 0.2473
N696 0.1268
N697 0.1243
N700 0.2473
N704 0.1249
N705 0.1243
N708 0.2473
N712 0.2301
N713 0.1243
N717 0.2473
N721 0.2301
N722 0.1243
N727 0.2473
N731 0.2301
N732 0.2186
N733 0.1649
N734 0.1164
N735 0.1263
N736 0.1999
N737 0.0686
N738 0.1263
N739 0.1999
N740 0.0686
N741 0.1263
N742 0.1999
N743 0.0686
N744 0.1263
N745 0.1999
N746 0.0686
N747 0.1243
N748 0.1997
N749 0.0674
N750 0.1243
N751 0.1997
N752 0.0674
N753 0.1243
N754 0.1997
N755 0.0674
N756 0.1243
N757 0.1739
N758 0.1997
N759 0.1997
N760 0.0674
N761 0.085
N762 0.085
N763 0.0569
N764 0.0869
N765 0.0869
N766 0.0584
N769 0.221
N770 0.221
N771 0.221
N772 0.221
N773 0.2332
N777 0.2206
N778 0.2372
N781 0.2206
N782 0.2438
N785 0.2206
N786 0.2462
N787 0.2206
N788 0.2026
N789 0.1625
N790 0.1993
N791 0.1679
N792 0.1922
N793 0.1783
N794 0.202
N795 0.1819
N796 0.2274
N802 0.245
N803 0.2451
N804 0.2453
N805 0.2485
N806 0.2064
N807 0.1558
N808 0.204
N809 0.2038
N810 0.2034
N811 0.1781
N812 0.1753
N813 0.1253
N814 0.0862
N815 0.2265
N819 0.2254
N822 0.2248
N825 0.2448
N826 0.2487
N827 0.2487
N828 0.2486
N829 0.1781
N830 0.207
N831 0.1548
N832 0.2076
N833 0.1536
N834 0.208
N835 0.1529
N836 0.2042
N837 0.2128
N838 0.1774
N839 0.1776
N840 0.1781
N841 0.1743
N842 0.2448
N843 0.2448
N844 0.2448
N845 0.2487
N846 0.2128
N847 0.1774
N848 0.1776
N849 0.2243
N851 0.2042
N852 0.2042
N853 0.2042
N854 0.2122
N855 0.2128
N856 0.1774
N857 0.1776
N858 0.2243
N859 0.2487
N860 0.2487
N861 0.2487
N862 0.2122
N867 0.2121
N868 0.2121
N869 0.2121
N870 0.2122
N871 0.2121
N872 0.2121
N873 0.2121
N875 0.2121
N876 0.2121
N877 0.2121


activity factors of the outputs: 
N388 0.1094
N389 0.1094
N390 0.1094
N391 0.1875
N418 0.0586
N419 0.0517
N420 0.1094
N421 0.1094
N422 0.1094
N423 0.2344
N446 0.0078
N447 0.1094
N448 0.0154
N449 0.0078
N450 0.2344
N767 0.2472
N768 0.2472
N850 0.1781
N863 0.2128
N864 0.1774
N865 0.1776
N866 0.2243
N874 0.2122
N878 0.2121
N879 0.2121
N880 0.2121


(base) bhaavanaa@bhaavanaa:~/VLSI_lab/DA2$*/
